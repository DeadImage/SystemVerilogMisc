package essentials;
	localparam LENGTH = 256;
endpackage